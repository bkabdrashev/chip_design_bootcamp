localparam RS =  546748 ;
