package alu_defines;
  localparam ALU_OP_END  = 3; 
  localparam ALU_OP_ADD  = 4'b0000; 
  localparam ALU_OP_SLL  = 4'b0001; 
  localparam ALU_OP_SLT  = 4'b0010; 
  localparam ALU_OP_SLTU = 4'b0011; 
  localparam ALU_OP_XOR  = 4'b0100; 
  localparam ALU_OP_SRL  = 4'b0101; 
  localparam ALU_OP_OR   = 4'b0110; 
  localparam ALU_OP_AND  = 4'b0111; 
  localparam ALU_OP_ANDN = 4'b1111; 
  localparam ALU_OP_LHS  = 4'b1010; 
  localparam ALU_OP_RHS  = 4'b1011; 
  localparam ALU_OP_SUB  = 4'b1000; 
  localparam ALU_OP_SRA  = 4'b1101; 
endpackage

