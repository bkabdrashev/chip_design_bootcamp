package com_defines;
  localparam COM_OP_END = 2; 
  localparam COM_OP_ONE = 3'b010; 
  localparam COM_OP_EQ  = 3'b000; 
  localparam COM_OP_NE  = 3'b001; 
  localparam COM_OP_LT  = 3'b100; 
  localparam COM_OP_GE  = 3'b101; 
  localparam COM_OP_LTU = 3'b110; 
  localparam COM_OP_GEU = 3'b111; 
endpackage

