localparam RS =  579211 ;
