localparam RS =  599521 ;
