module miniRV (
  input logic reset,
  input logic clk,
  input logic rom_wen,
  input logic rom_reset,
  input logic [31:0] rom_wdata,
  input logic [31:0] rom_addr,
  output logic [31:0] regs_out [0:15],
  output logic [31:0] pc,
  output logic [31:0] inst
);

  logic [4:0] dec_rd;
  logic [4:0] dec_rs1;
  logic [4:0] dec_rs2;
  logic [31:0] dec_imm;
  logic        dec_wen;
  logic [6:0]  dec_opcode;
  logic [2:0]  dec_funct3;

  logic is_pc_jump;
  logic [31:0]  pc_addr;

  logic [31:0] rdata1;
  logic [31:0] rdata2;
  logic [31:0] alu_res;

  logic [31:0] rom_addr_or_pc;

  logic [31:0] wdata;

  logic        ram_wen;
  logic [31:0] ram_addr;
  logic [31:0] ram_wdata;
  logic [31:0] ram_rdata;
  logic [3:0]  ram_wstrb;

  logic        vga_wen;
  logic [31:0] vga_addr;
  logic [31:0] vga_wdata;
  logic [31:0] vga_rdata;
  logic [3:0]  vga_wstrb;

  pc u_pc(
    .clk(clk),
    .reset(reset),
    .in_addr(pc_addr),
    .is_addr(is_pc_jump),
    .out_addr(pc)
  );

  ram64k #(.HEXFILE("vga2.hex")) ram(.clk(clk), .reset(reset),     .wen(ram_wen), .wdata(ram_wdata), .wstrb(ram_wstrb), .addr(ram_addr),       .read_data(ram_rdata));
  ram64k #(.HEXFILE("vga2.hex")) rom(.clk(clk), .reset(rom_reset), .wen(rom_wen), .wdata(rom_wdata), .wstrb(4'b1111),   .addr(rom_addr_or_pc), .read_data(inst));
  ram64k         #(.HEXFILE("")) vga(.clk(clk), .reset(reset),     .wen(vga_wen), .wdata(vga_wdata), .wstrb(vga_wstrb), .addr(vga_addr),       .read_data(vga_rdata));

  dec u_dec(
    .inst(inst),

    .rd(dec_rd),
    .rs1(dec_rs1),
    .rs2(dec_rs2),
    .imm(dec_imm),
    .wen(dec_wen),
    .opcode(dec_opcode),
    .funct3(dec_funct3)
  );

  alu u_alu(
    .opcode(dec_opcode),
    .rdata1(rdata1),
    .rdata2(rdata2),
    .imm(dec_imm),

    .rout(alu_res)
  );

  rf u_rf(
    .clk(clk),
    .reset(reset),
    .wen(dec_wen),
    .rd(dec_rd),
    .wdata(wdata),
    .rs1(dec_rs1),
    .rs2(dec_rs2),

    .rdata1(rdata1),
    .rdata2(rdata2),
    .regs_out(regs_out)
  );

  always_comb begin
    if (rom_wen) begin
      rom_addr_or_pc = rom_addr;

      ram_wen = 0;
      ram_addr = 0;
      ram_wdata = 0;
      ram_wstrb = 4'b0000;

      vga_wen = 0;
      vga_addr = 0;
      vga_wdata = 0;
      vga_wstrb = 0;

      wdata = 0;
      pc_addr = 0;
      is_pc_jump = 0;

    end else begin
      rom_addr_or_pc = pc;
      if (dec_opcode == 7'b0010011) begin
        // ADDI
        ram_wen = 0;
        ram_addr = 0;
        ram_wdata = 0;
        ram_wstrb = 4'b0000;

        vga_wen = 0;
        vga_addr = 0;
        vga_wdata = 0;
        vga_wstrb = 0;

        wdata = alu_res;
        pc_addr = 0;
        is_pc_jump = 0;
      end else if (dec_opcode == 7'b1100111) begin
        // JALR
        ram_wen = 0;
        ram_addr = 0;
        ram_wdata = 0;
        ram_wstrb = 0;

        vga_wen = 0;
        vga_addr = 0;
        vga_wdata = 0;
        vga_wstrb = 0;

        wdata = pc+4;
        pc_addr = (rdata1 + dec_imm) & ~3;
        is_pc_jump = 1;
      end else if (dec_opcode == 7'b0110011) begin
        // ADD
        ram_wen = 0;
        ram_addr = 0;
        ram_wdata = 0;
        ram_wstrb = 4'b0000;

        vga_wen = 0;
        vga_addr = 0;
        vga_wdata = 0;
        vga_wstrb = 0;

        wdata = alu_res;
        pc_addr = 0;
        is_pc_jump = 0;
      end else if (dec_opcode == 7'b0110111) begin
        // LUI
        ram_wen = 0;
        ram_addr = 0;
        ram_wdata = 0;
        ram_wstrb = 4'b0000;

        vga_wen = 0;
        vga_addr = 0;
        vga_wdata = 0;
        vga_wstrb = 0;

        wdata = dec_imm;
        pc_addr = 0;
        is_pc_jump = 0;
      end else if (dec_opcode == 7'b0000011 && dec_funct3 == 3'b010) begin
        // LW
        ram_wen = 0;
        ram_wdata = 0;
        ram_wstrb = 4'b0000;

        vga_wen = 0;
        vga_wdata = 0;
        vga_wstrb = 0;

        if (rdata1 + dec_imm < 'h2000_0000) begin
          ram_addr = rdata1 + dec_imm;
          vga_addr = 0;
          wdata = ram_rdata;
        end else begin
          ram_addr = 0;
          vga_addr = rdata1 + dec_imm - 'h2000_0000;
          wdata = vga_rdata;
        end

        pc_addr = 0;
        is_pc_jump = 0;
      end else if (dec_opcode == 7'b0000011 && dec_funct3 == 3'b100) begin
        // LBU
        ram_wen = 0;
        ram_wdata = 0;
        ram_wstrb = 0;

        vga_wen = 0;
        vga_wdata = 0;
        vga_wstrb = 0;

        if (rdata1 + dec_imm < 'h2000_0000) begin
          ram_addr = rdata1 + dec_imm;
          vga_addr = 0;
          wdata = ram_rdata & 32'hff;
        end else begin
          ram_addr = 0;
          vga_addr = rdata1 + dec_imm - 'h2000_0000;
          wdata = vga_rdata & 32'hff;
        end

        pc_addr = 0;
        is_pc_jump = 0;
      end else if (dec_opcode == 7'b0100011 && dec_funct3 == 3'b010) begin
        // SW
        if (rdata1 + dec_imm < 'h2000_0000) begin
          ram_wen = 1;
          ram_addr = rdata1 + dec_imm;
          ram_wdata = rdata2;
          ram_wstrb = 4'b1111;

          vga_wen = 0;
          vga_addr = 0;
          vga_wdata = 0;
          vga_wstrb = 0;
        end else begin
          ram_wen = 0;
          ram_addr = 0;
          ram_wdata = 0;
          ram_wstrb = 0;

          vga_wen = 1;
          vga_addr = rdata1 + dec_imm - 'h2000_0000;
          vga_wdata = rdata2;
          vga_wstrb = 4'b1111;
        end

        wdata = 0;
        pc_addr = 0;
        is_pc_jump = 0;
      end else if (dec_opcode == 7'b0100011 && dec_funct3 == 3'b000) begin
        // SB
        if (rdata1 + dec_imm < 'h2000_0000) begin
          ram_wen = 1;
          ram_addr = rdata1 + dec_imm;
          ram_wdata = rdata2 & 32'hff;
          ram_wstrb = 4'b0001;

          vga_wen = 0;
          vga_addr = 0;
          vga_wdata = 0;
          vga_wstrb = 0;
        end else begin
          ram_wen = 0;
          ram_addr = 0;
          ram_wdata = 0;
          ram_wstrb = 0;

          vga_wen = 1;
          vga_addr = rdata1 + dec_imm - 'h2000_0000;
          vga_wdata = rdata2 & 32'hff;
          vga_wstrb = 4'b0001;
        end

        wdata = 0;
        pc_addr = 0;
        is_pc_jump = 0;
      end else begin
        // NOT IMPLEMENTED
        ram_wen = 0;
        ram_addr = 0;
        ram_wdata = 0;
        ram_wstrb = 4'b0000;

        vga_wen = 0;
        vga_addr = 0;
        vga_wdata = 0;
        vga_wstrb = 0;

        wdata = 0;
        pc_addr = 0;
        wdata = 0;
        is_pc_jump = 0;
      end
    end
  end

endmodule;


