localparam RS =  574967 ;
