localparam RS =  540432 ;
