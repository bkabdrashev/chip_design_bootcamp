localparam REG_W_END = 31;
localparam REG_A_END = 4;
